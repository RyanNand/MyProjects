// Create the interface that will communicate with the DUT
interface dut_if;

  // Create ports that the DUT will utilize
  logic clock, reset;
  logic cmd;
  logic [7:0] addr;
  logic [7:0] data;

endinterface

// Create the DUT or the device to be tested
module dut(dut_if dif);

  // Import in the UVM base class library
    // We are using "'uvm_info()" for reporting in the procedural block below
  import uvm_pkg::*;

  // Create a procedural block for reporting and your arbitrary design
    // Will trigger on the positive edge of clock provided through the interface
  always @(posedge dif.clock) begin
    // Report the values received from the interface
	  // In SystemVerilog, "$sformatf" is a system task that type casts data into a string format
	  // In SystemVerilog, "%b" is a binary value and "%d" is a decimal value
    `uvm_info("", $sformatf("DUT received cmd=%b, addr=%d, data=%d",
                            dif.cmd, dif.addr, dif.data), UVM_MEDIUM)
  end
  
endmodule
